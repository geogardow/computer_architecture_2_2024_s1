module mem_output_manager();


endmodule