
module flags (
	source,
	probe);	

	output	[18:0]	source;
	input	[18:0]	probe;
endmodule
